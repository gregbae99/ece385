module FontDriver (input        [4:0]   In0,
						 output logic [143:0] Out0);
	always_comb
	begin
		unique case (In0)
			5'b00000: Out0 = 144'b000000000000000111111000001111111100001100001100001100001100001100001100001100001100001100001100001100001100001111111100000111111000000000000000; //0
			5'b00001: Out0 = 144'b000000000000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000000000000; //1
			5'b00010: Out0 = 144'b000000000000000111111000001111111100000000001100000000001100000111111100001111111000001100000000001100000000001111111100000111111000000000000000; //2
			5'b00011: Out0 = 144'b000000000000000111111000001111111100000000001100000000001100000111111100000111111100000000001100000000001100001111111100000111111000000000000000; //3
			5'b00100: Out0 = 144'b000000000000001100001100001100001100001100001100001100001100001111111100000111111100000000001100000000001100000000001100000000001100000000000000; //4
			5'b00101: Out0 = 144'b000000000000000111111000001111111100001100000000001100000000001111111000000111111100000000001100000000001100001111111100000111111000000000000000; //5
			5'b00110: Out0 = 144'b000000000000000111111000001111111100001100000000001100000000001111111000001111111100001100001100001100001100001111111100000111111000000000000000; //6
			5'b00111: Out0 = 144'b000000000000000111111000001111111100001100001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000000000; //7
			5'b01000: Out0 = 144'b000000000000000111111000001111111100001100001100001100001100001111111100001111111100001100001100001100001100001111111100000111111000000000000000; //8
			5'b01001: Out0 = 144'b000000000000000111111000001111111100001100001100001100001100001111111100001111111100000000001100000000001100001111111100000111111000000000000000; //9
			5'b10001: Out0 = 144'b000000000000000111111000001111111100001100001100001100001100001111111100001111111000001100000000001100000000001100000000001100000000000000000000; //P
			5'b10010: Out0 = 144'b000000000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001111111100000111111000000000000000; //L
			5'b10011: Out0 = 144'b000000000000000111111000001111111100001100001100001100001100001111111100001111111100001100001100001100001100001100001100001100001100000000000000; //A
			5'b10100: Out0 = 144'b000000000000001100001100001100001100001100001100001100001100001111111100000111111000000001100000000001100000000001100000000001100000000000000000; //Y
			5'b10101: Out0 = 144'b000000000000000111111000001111111100001100000000001100000000001111111100001111111100001100000000001100000000001111111100000111111000000000000000; //E
			5'b10110: Out0 = 144'b000000000000000111111000001111111100001100001100001100001100001111111100001111111100001100011000001100001100001100001100001100001100000000000000; //R
			5'b10111: Out0 = 144'b000000000000000111111000001111111100001100000000001100000000001100111100001100111100001100001100001100001100001111111100000111111000000000000000; //G
			5'b11000: Out0 = 144'b000000000000000110011000001111111100001101101100001101101100001101101100001101101100001101101100001101101100001101101100001101101100000000000000; //M
			5'b11001: Out0 = 144'b000000000000001100001100001100001100001100001100001100001100000110011000000110011000000110011000000011110000000011110000000001100000000000000000; //V
			5'b11010: Out0 = 144'b000000000000001101101100001101101100001101101100001101101100001101101100001101101100001101101100001101101100001111111100000110011000000000000000; //W
			5'b11011: Out0 = 144'b000000000000001100001100001100001100001110001100001111001100001101101100001101101100001100111100001100011100001100001100001100001100000000000000; //N
			5'b11100: Out0 = 144'b000000000000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000000000000000001100000000001100000000000000000; //!
			5'b11101: Out0 = 144'b000000000000011111111110011111111110011111111110011111111110011111111110011111111110011111111110011111111110011111111110011111111110000000000000; //Block
			default: Out0 = 144'b0; //Empty
		endcase
	end
endmodule
